library verilog;
use verilog.vl_types.all;
entity MeioSomador_vlg_vec_tst is
end MeioSomador_vlg_vec_tst;
