library verilog;
use verilog.vl_types.all;
entity MeioSomador_vlg_check_tst is
    port(
        s               : in     vl_logic;
        Ts              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MeioSomador_vlg_check_tst;
